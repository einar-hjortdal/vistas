module main

const plausible_gzip = ['.html', '.css', '.js', '.json', '.xml', '.md']
const gzip_extension = '.gz'
