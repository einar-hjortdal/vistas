module main

const plausible_gzip = ['.html', '.css', '.js', '.json', '.xml', '.md', '.txt']
const gzip_extension = '.gz'
