module main

// import net.http

fn parse_authorization_header(authorization string) {
}

// fn validate_signature() {
//	authorization := ctx.get_header(http.CommonHeader.authorization) or { return error }
// parse_authorization_header(authorization) or { return error }
// }
